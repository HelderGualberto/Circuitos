library verilog;
use verilog.vl_types.all;
entity halfSubtractor_vlg_vec_tst is
end halfSubtractor_vlg_vec_tst;
