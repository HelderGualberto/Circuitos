library verilog;
use verilog.vl_types.all;
entity adder7b_vlg_vec_tst is
end adder7b_vlg_vec_tst;
