library verilog;
use verilog.vl_types.all;
entity UnidadedeControle_vlg_vec_tst is
end UnidadedeControle_vlg_vec_tst;
