library verilog;
use verilog.vl_types.all;
entity Mux5to1_vlg_vec_tst is
end Mux5to1_vlg_vec_tst;
