library verilog;
use verilog.vl_types.all;
entity andFunction_vlg_vec_tst is
end andFunction_vlg_vec_tst;
