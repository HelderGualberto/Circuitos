library verilog;
use verilog.vl_types.all;
entity comp2_vlg_vec_tst is
end comp2_vlg_vec_tst;
