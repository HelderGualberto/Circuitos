library verilog;
use verilog.vl_types.all;
entity Integracao_vlg_vec_tst is
end Integracao_vlg_vec_tst;
