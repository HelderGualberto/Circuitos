library verilog;
use verilog.vl_types.all;
entity orFunction_vlg_vec_tst is
end orFunction_vlg_vec_tst;
