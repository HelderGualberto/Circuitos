library verilog;
use verilog.vl_types.all;
entity dataFlux_vlg_vec_tst is
end dataFlux_vlg_vec_tst;
