library verilog;
use verilog.vl_types.all;
entity orFunction_vlg_check_tst is
    port(
        S               : in     vl_logic_vector(0 to 6);
        sampler_rx      : in     vl_logic
    );
end orFunction_vlg_check_tst;
