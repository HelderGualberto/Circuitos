library verilog;
use verilog.vl_types.all;
entity UFA_vlg_vec_tst is
end UFA_vlg_vec_tst;
