library verilog;
use verilog.vl_types.all;
entity teste is
    port(
        CLKFD           : out    vl_logic;
        CLKUC           : in     vl_logic
    );
end teste;
