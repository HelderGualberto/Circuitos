library verilog;
use verilog.vl_types.all;
entity register7b_vlg_vec_tst is
end register7b_vlg_vec_tst;
