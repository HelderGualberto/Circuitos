library verilog;
use verilog.vl_types.all;
entity mux8bits_vlg_vec_tst is
end mux8bits_vlg_vec_tst;
