library verilog;
use verilog.vl_types.all;
entity FluxoDeDados_vlg_vec_tst is
end FluxoDeDados_vlg_vec_tst;
