library verilog;
use verilog.vl_types.all;
entity subtractor7b_vlg_vec_tst is
end subtractor7b_vlg_vec_tst;
